magic
tech sky130A
timestamp 1628502354
<< nwell >>
rect 319 256 473 258
rect -257 243 473 256
rect -257 172 475 243
rect -256 125 475 172
rect 36 115 475 125
rect 251 114 475 115
rect -76 -277 74 -276
rect -115 -278 121 -277
rect -118 -279 121 -278
rect 290 -279 475 114
rect -118 -414 475 -279
rect -118 -423 474 -414
rect -115 -424 86 -423
rect -76 -425 74 -424
rect 263 -425 474 -423
<< nmos >>
rect -23 -117 27 -74
<< pmos >>
rect -23 -402 27 -301
<< ndiff >>
rect -237 -41 -184 -8
rect -184 -364 -182 -42
rect -82 -76 -23 -74
rect -83 -83 -23 -76
rect -83 -107 -79 -83
rect -50 -107 -23 -83
rect -83 -117 -23 -107
rect 27 -85 81 -74
rect 27 -109 46 -85
rect 75 -109 81 -85
rect 27 -117 81 -109
rect -253 -365 -182 -364
<< pdiff >>
rect -100 -308 -23 -301
rect -100 -332 -88 -308
rect -59 -332 -23 -308
rect -100 -364 -23 -332
rect -100 -388 -86 -364
rect -57 -388 -23 -364
rect -100 -401 -23 -388
rect -51 -402 -23 -401
rect 27 -307 102 -301
rect 27 -331 63 -307
rect 92 -331 102 -307
rect 27 -363 102 -331
rect 27 -387 62 -363
rect 91 -387 102 -363
rect 27 -401 102 -387
rect 27 -402 54 -401
rect 37 -403 54 -402
<< ndiffc >>
rect -240 14 -194 56
rect 49 39 84 65
rect 156 61 180 81
rect -242 -162 -196 -110
rect -237 -349 -191 -307
rect 49 -24 83 3
rect 159 -25 182 -2
rect -79 -107 -50 -83
rect 46 -109 75 -85
rect -89 -481 -60 -460
rect -85 -574 -56 -553
<< pdiffc >>
rect -88 -332 -59 -308
rect -86 -388 -57 -364
rect 63 -331 92 -307
rect 62 -387 91 -363
<< nsubdiff >>
rect -78 168 -21 174
rect -78 149 -63 168
rect -39 149 -21 168
rect -78 143 -21 149
<< nsubdiffcont >>
rect -63 149 -39 168
<< poly >>
rect -23 -30 27 -12
rect -23 -50 -11 -30
rect 14 -50 27 -30
rect -23 -74 27 -50
rect -23 -133 27 -117
rect -23 -227 27 -204
rect -23 -251 -11 -227
rect 18 -251 27 -227
rect -23 -301 27 -251
rect -23 -416 27 -402
<< polycont >>
rect -11 -50 14 -30
rect -11 -251 18 -227
<< ndiffres >>
rect -253 56 -182 83
rect 149 81 188 91
rect -253 14 -240 56
rect -194 14 -182 56
rect -253 -8 -182 14
rect -253 -41 -237 -8
rect -184 -41 -182 -8
rect 38 65 97 75
rect 38 39 49 65
rect 84 39 97 65
rect 149 61 156 81
rect 180 61 188 81
rect 149 51 188 61
rect 38 3 97 39
rect -253 -42 -182 -41
rect -253 -110 -184 -42
rect -253 -162 -242 -110
rect -196 -162 -184 -110
rect -253 -307 -184 -162
rect -253 -349 -237 -307
rect -191 -349 -184 -307
rect -253 -364 -184 -349
rect 38 -24 49 3
rect 83 -7 97 3
rect 148 -2 188 51
rect 83 -24 96 -7
rect 38 -30 96 -24
rect 148 -25 159 -2
rect 182 -25 188 -2
rect 148 -33 188 -25
rect -99 -460 -49 -451
rect -99 -481 -89 -460
rect -60 -481 -49 -460
rect -99 -553 -49 -481
rect -99 -574 -85 -553
rect -56 -574 -49 -553
rect -99 -579 -49 -574
<< locali >>
rect -255 193 175 194
rect -256 174 175 193
rect -255 168 175 174
rect -255 161 -63 168
rect -255 135 -232 161
rect -200 149 -63 161
rect -39 154 175 168
rect -39 149 133 154
rect -200 135 133 149
rect -255 128 133 135
rect 167 128 175 154
rect -255 115 175 128
rect -250 67 -188 115
rect 150 91 175 115
rect 150 89 188 91
rect 149 81 188 89
rect -66 70 -22 80
rect 43 70 93 74
rect -251 56 -189 67
rect -251 14 -240 56
rect -194 14 -189 56
rect -66 66 93 70
rect -66 39 -57 66
rect -32 65 93 66
rect -32 39 49 65
rect 84 58 93 65
rect 149 61 156 81
rect 180 61 188 81
rect 84 39 132 58
rect 149 51 188 61
rect -66 38 132 39
rect -66 28 -22 38
rect 43 36 132 38
rect 43 29 98 36
rect -251 1 -189 14
rect 49 11 89 12
rect 42 3 97 11
rect -20 -23 22 -20
rect -144 -30 22 -23
rect 42 -24 49 3
rect 83 -24 97 3
rect 42 -29 97 -24
rect -144 -50 -11 -30
rect 14 -50 22 -30
rect 43 -31 97 -29
rect 115 10 132 36
rect 115 9 133 10
rect 115 7 149 9
rect 115 -2 188 7
rect 115 -25 159 -2
rect 182 -25 188 -2
rect 43 -32 74 -31
rect -144 -55 22 -50
rect -144 -56 21 -55
rect -252 -110 -185 -103
rect -252 -162 -242 -110
rect -196 -126 -185 -110
rect -144 -126 -117 -56
rect 53 -74 74 -32
rect 115 -34 188 -25
rect -82 -75 -45 -74
rect -83 -83 -45 -75
rect -83 -107 -79 -83
rect -50 -107 -45 -83
rect -83 -117 -45 -107
rect 42 -85 80 -74
rect 42 -109 46 -85
rect 75 -109 80 -85
rect 42 -117 80 -109
rect -196 -156 -117 -126
rect -196 -157 -118 -156
rect -196 -162 -185 -157
rect -252 -168 -185 -162
rect -81 -218 -45 -117
rect -81 -227 46 -218
rect -81 -251 -11 -227
rect 18 -251 46 -227
rect -81 -260 46 -251
rect 148 -279 182 -34
rect -246 -292 -184 -290
rect -248 -307 -184 -292
rect -248 -349 -237 -307
rect -191 -349 -184 -307
rect -248 -358 -184 -349
rect -99 -308 -47 -301
rect -99 -332 -88 -308
rect -59 -332 -47 -308
rect -234 -605 -187 -358
rect -99 -364 -47 -332
rect -99 -388 -86 -364
rect -57 -388 -47 -364
rect -99 -400 -47 -388
rect 50 -307 102 -301
rect 148 -307 183 -279
rect 50 -331 63 -307
rect 92 -331 183 -307
rect 50 -336 183 -331
rect 50 -363 102 -336
rect 50 -387 62 -363
rect 91 -387 102 -363
rect 50 -400 102 -387
rect -84 -451 -61 -400
rect -98 -460 -52 -451
rect -98 -481 -89 -460
rect -60 -481 -52 -460
rect -98 -494 -52 -481
rect -97 -548 -50 -545
rect -99 -553 -50 -548
rect -99 -574 -85 -553
rect -56 -564 -50 -553
rect -56 -574 -49 -564
rect -99 -605 -49 -574
rect -234 -617 -49 -605
rect -234 -636 -222 -617
rect -190 -618 -49 -617
rect -190 -636 -91 -618
rect -234 -638 -91 -636
rect -54 -638 -49 -618
rect -234 -645 -49 -638
<< viali >>
rect -232 135 -200 161
rect 133 128 167 154
rect -57 39 -32 66
rect -222 -636 -190 -617
rect -91 -638 -54 -618
<< metal1 >>
rect -254 173 173 193
rect -256 161 175 173
rect -256 135 -232 161
rect -200 154 175 161
rect -200 135 133 154
rect -256 128 133 135
rect 167 128 175 154
rect -256 115 175 128
rect -65 66 -25 78
rect -65 39 -57 66
rect -32 39 -25 66
rect -65 29 -25 39
rect -234 -617 -49 -607
rect -234 -636 -222 -617
rect -190 -618 -49 -617
rect -190 -636 -91 -618
rect -234 -638 -91 -636
rect -54 -638 -49 -618
rect -234 -646 -49 -638
<< labels >>
rlabel viali -230 139 -209 151 1 vdd
rlabel viali -54 41 -40 58 1 out
rlabel ndiffc -238 -155 -201 -120 1 in
rlabel metal1 -222 -637 -194 -619 1 gnd
<< end >>
