* SPICE3 file created from spamp.ext - technology: sky130A

.option scale=10000u

X0 a_27_n117# out SUB sky130_fd_pr__res_generic_nd w=34 l=36
X1 vdd a_n237_n41# SUB sky130_fd_pr__res_generic_nd w=46 l=22
X2 out a_n83_n117# a_n100_n401# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=50
X3 vdd out SUB sky130_fd_pr__res_generic_nd w=22 l=63
X4 a_n100_n401# gnd SUB sky130_fd_pr__res_generic_nd w=27 l=72
X5 a_27_n117# in a_n83_n117# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=42 l=50
C0 vdd SUB 4.11fF
