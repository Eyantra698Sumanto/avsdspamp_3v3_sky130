magic
tech sky130A
timestamp 1629117458
<< nwell >>
rect -2673 6125 2341 7034
rect -185 200 86 6125
rect -286 -136 347 200
<< nmos >>
rect -1344 207 -1244 307
<< pmos >>
rect -27 -97 73 3
<< ndiff >>
rect -1544 282 -1344 307
rect -1544 228 -1536 282
rect -1482 228 -1344 282
rect -1544 207 -1344 228
rect -1244 280 -1044 307
rect -1244 227 -1118 280
rect -1064 227 -1044 280
rect -1244 207 -1044 227
<< pdiff >>
rect -123 -19 -27 3
rect -123 -71 -116 -19
rect -75 -71 -27 -19
rect -123 -97 -27 -71
rect 73 -21 177 3
rect 73 -73 122 -21
rect 163 -73 177 -21
rect 73 -97 177 -73
<< ndiffc >>
rect -1536 228 -1482 282
rect -1118 227 -1064 280
<< pdiffc >>
rect -116 -71 -75 -19
rect 122 -73 163 -21
<< nsubdiff >>
rect -545 6554 832 6592
rect -545 6403 -160 6554
rect 49 6403 832 6554
rect -545 6321 832 6403
<< nsubdiffcont >>
rect -160 6403 49 6554
<< poly >>
rect -1344 307 -1244 385
rect -1344 -28 -1244 207
rect -27 3 73 42
rect -1344 -75 -1313 -28
rect -1271 -75 -1244 -28
rect -1344 -115 -1244 -75
rect -27 -389 73 -97
rect -27 -441 10 -389
rect 49 -441 73 -389
rect -27 -458 73 -441
<< polycont >>
rect -1313 -75 -1271 -28
rect 10 -441 49 -389
<< xpolycontact >>
rect -1153 5717 -973 6081
rect -2355 4764 -2160 5124
rect 1178 5065 1341 5421
rect -1175 383 -995 747
rect 2039 4956 2208 5310
rect -2355 -482 -2160 -122
rect 1171 -163 1356 207
rect 2017 -496 2186 -142
<< xpolyres >>
rect -2306 -122 -2271 4764
rect -1092 747 -1057 5717
rect 1261 207 1296 5065
rect 2122 -142 2157 4956
<< locali >>
rect -2086 6668 1949 6737
rect -2086 6358 -1972 6668
rect -1581 6554 1482 6668
rect -1581 6403 -160 6554
rect 49 6403 1482 6554
rect -1581 6358 1482 6403
rect -2086 6352 1482 6358
rect 1855 6352 1949 6668
rect -2086 6295 1949 6352
rect -1157 6081 -968 6295
rect -1157 6067 -1153 6081
rect -1159 5868 -1153 6067
rect -2711 5822 -1486 5828
rect -3412 5664 -1486 5822
rect -973 6067 -968 6081
rect -973 5868 -966 6067
rect -3412 5361 -3311 5664
rect -2982 5645 -1486 5664
rect -2982 5361 -1909 5645
rect -3412 5342 -1909 5361
rect -1580 5342 -1486 5645
rect 1614 5462 1880 6295
rect -3412 5222 -1486 5342
rect 671 5264 933 5276
rect -3412 5216 -2187 5222
rect -2364 5124 -2187 5216
rect 671 5151 1178 5264
rect -2364 4925 -2355 5124
rect -2160 4917 -1542 4943
rect -2160 4764 -1478 4917
rect -2344 4752 -1478 4764
rect -1657 282 -1478 4752
rect -598 1168 -450 1217
rect -598 1112 -548 1168
rect -505 1112 -450 1168
rect -598 655 -450 1112
rect 671 655 933 5151
rect 1614 5329 2183 5462
rect 1614 5317 1880 5329
rect 2031 5310 2176 5329
rect 2031 5127 2039 5310
rect -830 513 945 655
rect -1657 228 -1536 282
rect -1482 228 -1478 282
rect -1657 168 -1478 228
rect -1141 280 -1037 383
rect -1141 227 -1118 280
rect -1064 227 -1037 280
rect -1141 211 -1037 227
rect -1141 177 -1040 211
rect -1321 9 -68 10
rect -1365 2 -68 9
rect 108 2 1171 12
rect -1365 -19 -55 2
rect -1365 -28 -116 -19
rect -1365 -75 -1313 -28
rect -1271 -71 -116 -28
rect -75 -71 -55 -19
rect -1271 -75 -55 -71
rect -1365 -97 -55 -75
rect 107 -21 1171 2
rect 107 -73 122 -21
rect 163 -73 1171 -21
rect 107 -97 1171 -73
rect -1365 -99 -68 -97
rect 108 -109 1171 -97
rect -2466 -454 -2355 -360
rect -2160 -365 -2138 -360
rect -2160 -368 33 -365
rect -2160 -389 2017 -368
rect -2160 -441 10 -389
rect 49 -441 2017 -389
rect -2160 -451 2017 -441
rect -2160 -454 79 -451
rect -30 -740 79 -454
rect 2186 -451 2227 -368
rect -30 -786 2 -740
rect 57 -786 79 -740
rect -30 -805 79 -786
<< viali >>
rect -1972 6358 -1581 6668
rect 1482 6352 1855 6668
rect -3311 5361 -2982 5664
rect -1909 5342 -1580 5645
rect -548 1112 -505 1168
rect 2 -786 57 -740
<< metal1 >>
rect -2086 6668 1949 6737
rect -2086 6358 -1972 6668
rect -1581 6358 1482 6668
rect -2086 6352 1482 6358
rect 1855 6352 1949 6668
rect -2086 6295 1949 6352
rect -2711 5822 -1486 5828
rect -3412 5664 -1486 5822
rect -3412 5361 -3311 5664
rect -2982 5645 -1486 5664
rect -2982 5361 -1909 5645
rect -3412 5342 -1909 5361
rect -1580 5342 -1486 5645
rect -3412 5222 -1486 5342
rect -3412 5216 -2187 5222
rect -598 1168 -462 1211
rect -598 1112 -548 1168
rect -505 1112 -462 1168
rect -598 1075 -462 1112
rect -50 -740 109 -714
rect -50 -786 2 -740
rect 57 -786 109 -740
rect -50 -811 109 -786
<< labels >>
rlabel metal1 3 -786 58 -740 1 vin
rlabel viali -548 1112 -505 1168 1 vout
rlabel metal1 -255 6390 143 6617 1 vdd
rlabel metal1 -2648 5354 -2269 5582 1 gnd
<< end >>
