magic
tech sky130A
timestamp 1629117458
<< labels >>
rlabel metal1 3 -786 58 -740 1 vin
rlabel viali -548 1112 -505 1168 1 vout
rlabel metal1 -255 6390 143 6617 1 vdd
rlabel metal1 -2648 5354 -2269 5582 1 gnd
<< end >>
