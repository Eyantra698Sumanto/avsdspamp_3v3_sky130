* SPICE3 file created from /home/sumanto/Desktop/layout/spamp.ext - technology: sky130A
.lib "sky130_fd_pr/models/sky130.lib.spice" tt
* SPICE3 file created from /home/sumanto/Desktop/layout/spamp.ext - technology: sky130A

X0 a_27_n117# out SUB sky130_fd_pr__res_generic_nd w=34 l=36
X1 vdd a_n237_n41# SUB sky130_fd_pr__res_generic_nd w=46 l=22
X2 out a_n83_n117# a_n100_n401# vdd sky130_fd_pr__pfet_01v8  w=100 l=50
X3 vdd out SUB sky130_fd_pr__res_generic_nd w=22 l=63
*vo out vdd 0; Current Gain Vs Collector Current 
X4 a_n100_n401# gnd SUB sky130_fd_pr__res_generic_nd w=27 l=72
X5 a_27_n117# in a_n83_n117# SUB sky130_fd_pr__nfet_01v8  w=42 l=50
C0 vdd SUB 4.11fF

v2 vdd gnd dc 1.8; Supply for Transient, AC analysis 
*v2 vdd gnd 0 pwl (0 0 100m 3); Variation of supply analysis 
v1 in gnd sine(0 10m 100 0 0); for Transient analysis 
* v1 in gnd 1; Variation of supply analysis 
* I1 in gnd 1; Current Gain Vs Collector Current
* v1 in gnd dc 0 ac 10m; for AC analysis 
.tran 10e-06 100e-03 0e-03; for Transient analysis, supply 
variation analysis
*.temp 50;
.control;
run;
print allv > plot_data_v.txt;
print alli > plot_data_i.txt;
*ac dec 100 1 100Meg; AC analysis 
*plot vdb(out)/vdb(in); AC analysis 
plot v(out) v(in); Transient Analysis 
*plot v(out) vs v(vdd); Variation of supply analysis 
*plot Vo#branch vs V2#branch; Current Gain Vs Collector Current 
.endc
.end